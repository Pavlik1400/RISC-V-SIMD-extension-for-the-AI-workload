// Default configuration for simc_v2 CNN_1 model
    // parameter INPUT_SIZE = 1024;
    // parameter MAX_INPUT_SIZE = INPUT_SIZE;

    // parameter PADDING = 4;  // (8 / 2)
    // parameter MAX_INPUT_CHANNELS = 128;
    // parameter KERNEL_LENGTH = 8;

// // Default configuration for radioml CNN_1 model
//     parameter INPUT_SIZE = 128;
//     parameter MAX_INPUT_SIZE = INPUT_SIZE;

//     parameter PADDING = 4;  // (8 / 2)
//     parameter MAX_INPUT_CHANNELS = 128;
//     parameter KERNEL_LENGTH = 8;

// Default configuration for radioml CNN_1 model small
    parameter INPUT_SIZE = 128;
    // parameter ACTUAL_MAX_INPUT_SIZE = 4096;
    parameter ACTUAL_MAX_INPUT_SIZE = 4352;
    // parameter ACTUAL_MAX_INPUT_SIZE = 8192;

    parameter PADDING = 4;  // (8 / 2)
    parameter MAX_INPUT_CHANNELS = 64;
    parameter KERNEL_LENGTH = 8;