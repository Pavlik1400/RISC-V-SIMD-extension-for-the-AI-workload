// Default configuration for simc_v2 CNN_1 model
    // parameter INPUT_SIZE = 1024;
    // parameter MAX_INPUT_SIZE = INPUT_SIZE;

    // parameter PADDING = 4;  // (8 / 2)
    // parameter MAX_INPUT_CHANNELS = 128;
    // parameter KERNEL_LENGTH = 8;

// Default configuration for radioml CNN_1 model
    parameter INPUT_SIZE = 128;
    parameter MAX_INPUT_SIZE = INPUT_SIZE;

    parameter PADDING = 4;  // (8 / 2)
    parameter MAX_INPUT_CHANNELS = 128;
    parameter KERNEL_LENGTH = 8;